library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity ParallelEnc is
port();
end ParallelEnc;

architecture Behavoral of ParallelEnc is
begin

end;