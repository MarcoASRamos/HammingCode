library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity ParallelDecod is
port();
end ParallelDecod;

architecture Behavoral of ParallelDecod is
begin

end;